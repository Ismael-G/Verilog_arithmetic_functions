lfkjak;li sdafsa
andslkjncj kasn


module verturned_staircase_tree_multiplication(
  
);

input logic product1 ;

input logic product2 ;

output logic result;

assign result = product1 * product2 ;


endmodule
