 /*
  * Ismael Garcia 
  * January 2021
  * weinberber multiplication is the use of a balanced tree in order to
  * compute multiplcation
  *
  */

module weinberber_multiplication(
  
);

input wire product1; 
input wire product2; 

output wire result ;


assign result = product1 * product2 ; 


endmodule
