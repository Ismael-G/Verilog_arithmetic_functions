 /* 
  * Ismael Garcia
  * January 2021
  * ldkjf
  * lksjadlkfj
  * lsdkjlf
  */
module wallace_tree(
  
);
input logic product1 ;
input logic product2 ;

output logic result;


assign result = product1 * product2 ;



endmodule
