/* 
  * Ismael Garcia
  * January 2021
  * Goldschmidt Division Algorithm implemented in system verilog
*/

module goldschmidt_division(
  
);

input logic dividend ;
input logic divisor ;

output logic quotient ; 


endmodule
