// test bench for the carry skip adder goes here
